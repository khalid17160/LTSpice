* E:\LTSpice\Upload\q1\q1,2_sch.asc
R1 0 N001 100
R2 N002 0 100
R3 N003 N002 70
R5 0 N002 220
R6 0 N003 150
V1 N001 0 10
.op
.backanno
.end
