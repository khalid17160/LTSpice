* E:\LTSpice\Upload_2_dead\clamper1\clamper.asc
V1 N001 0 PULSE(10 -10 10 0 0 10 20 100)
C1 vout N001 200�
D1 0 vout D
.model D D
.lib C:\Users\Khalid\Documents\LTspiceXVII\lib\cmp\standard.dio
.tran 100s
.backanno
.end
