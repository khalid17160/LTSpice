* E:\LTSpice\Upload\DiffernceAmp_sch.asc
XU1 N005 N001 P001 P002 N002 AD8066
R2 N001 N003 1k
V1 P001 0 20
V2 0 P002 12
R3 N002 0 10k
V3 N003 0 SINE(0 2 500)
R1 N002 N001 1K
V4 N004 0 SINE(0 5 500)
R4 N005 N004 1k
R5 N005 0 1k
.tran 10m
.lib ADI.lib
.backanno
.end
