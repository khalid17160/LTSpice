* E:\LTSpice\Upload\Draft1.asc
XU1 0 N001 P001 P002 N002 AD8066;
R1 N001 N003 2k;
R2 N002 N001 2K;
V1 P001 0 12;
V2 0 P002 12;
R3 N002 0 10k;
V3 N003 0 SINE(0 5 200);
.tran 10m;
.lib ADI.lib;
.backanno;
.end;
